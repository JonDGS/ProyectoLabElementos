* SPICE3 file created from nand.ext - technology: scmos

.option scale=0.3u

M1000 vout va VDD w_n24_n9# pfet w=18 l=3
+  ad=198 pd=58 as=342 ps=110
M1001 VDD vb vout w_n24_n9# pfet w=18 l=3
+  ad=0 pd=0 as=0 ps=0
M1002 vout vb a_n5_n39# Gnd nfet w=10 l=3
+  ad=110 pd=42 as=110 ps=42
M1003 a_n5_n39# va GND Gnd nfet w=10 l=3
+  ad=0 pd=0 as=80 ps=36
C0 w_n24_n9# Gnd 6.55fF
